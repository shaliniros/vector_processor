`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 26.04.2021 01:35:25
// Design Name: 
// Module Name: vector_proc
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`include "definitions.v"

module vector_proc();
     fetch      f1 ();
     decode     d1();
     execute    exe1();
     mem_access mem1();
     write_back wb1();
endmodule
